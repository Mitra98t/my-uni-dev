module hello (
    output z, 
    input a
);
    
    assign z = a;

endmodule